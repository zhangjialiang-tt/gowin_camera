parameter WIDTH_B = 16;
parameter DELAY = 5;
parameter WIDTH_A = 16;
