//Copyright (C)2014-2025 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.11.03 (64-bit)
//Part Number: GW2ANR-LV18QN88C8/I7
//Device: GW2ANR-18
//Device Version: C
//Created Time: Tue Sep 30 13:33:25 2025

module Gowin_pROM (dout, clk, oce, ce, reset, ad);

output [15:0] dout;
input clk;
input oce;
input ce;
input reset;
input [8:0] ad;

wire [15:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[15:0],dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({gw_gnd,ad[8:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 16;
defparam prom_inst_0.RESET_MODE = "ASYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h1B4B1A01190E18221714122E10520F060EC00D040C000B000A00090004E20304;
defparam prom_inst_0.INIT_RAM_01 = 256'h807F34013306319030012D6026102501241622A0214020031F781E881D101C07;
defparam prom_inst_0.INIT_RAM_02 = 256'hC746C63BC590C480C300B0558B008A0085088903880386038402830082FA8126;
defparam prom_inst_0.INIT_RAM_03 = 256'h410040429840970696B0950494009300920091009001B601EF90EE60ED04EC06;
defparam prom_inst_0.INIT_RAM_04 = 256'h6B086A08760069206820672066206500640063006200610060005F005E00435B;
defparam prom_inst_0.INIT_RAM_05 = 256'h0900FE014B0B49004815FE027F007E3C72F07600710870086F086E086D086C08;
defparam prom_inst_0.INIT_RAM_06 = 256'h15B01235FE010F04FE022320224020401F351E611C111700136B11100C100B11;
defparam prom_inst_0.INIT_RAM_07 = 256'h8205810880C1A21197659584943392CB9103906CFE02410F40903FB03E281031;
defparam prom_inst_0.INIT_RAM_08 = 256'hAB40A680A540A420A350FE022104FE018B108A3089B08815875086F0840A8308;
defparam prom_inst_0.INIT_RAM_09 = 256'h142713191213110D1009FE024C204B063D153C04B92BB701B638B464B346AE0C;
defparam prom_inst_0.INIT_RAM_0A = 256'h24F923F522EF21EA20E31FD91ECD1DBD1CA91B9D1A8F197D1869175316451537;
defparam prom_inst_0.INIT_RAM_0B = 256'h307C2F692E592D452C3B2B332A27291E28192714260FFE02C72BC620FE0025FF;
defparam prom_inst_0.INIT_RAM_0C = 256'hD710D6F0D340D232D1323BFF3AF939F338E937E236DA35CF34C033AE32983189;
defparam prom_inst_0.INIT_RAM_0D = 256'hBC24CA0AC90DC815C40CC30DC2149F40FE01D8D8EF3FEE00ED80DE86DD14D8DA;
defparam prom_inst_0.INIT_RAM_0E = 256'hBA00B900C100C000BF07CD00CC00CB00C700C600C500B815B716B625BE0BBD10;
defparam prom_inst_0.INIT_RAM_0F = 256'hD200D100D009B50EB40EB317B206B107B00BAF0EAE06AD05AC00AB01AA01BB00;
defparam prom_inst_0.INIT_RAM_10 = 256'hA180A977A877A777A677A500A400D500D400D30ADB00DA00D900D800D700D608;
defparam prom_inst_0.INIT_RAM_11 = 256'h4B014F004F00E9A0E890E7A0E690E390E277E180E077DD30DC25DF0DFE01A280;
defparam prom_inst_0.INIT_RAM_12 = 256'h4E024DB04C014E024D904C014E014D704C014E014D914C014E014D714C014F00;
defparam prom_inst_0.INIT_RAM_13 = 256'h4C014E024DF04C014E024DD04C014E024DAF4C014E024D6F4C014E024D8F4C01;
defparam prom_inst_0.INIT_RAM_14 = 256'h4DCE4C014E034DAE4C014E034D8E4C014E034D6E4C014E024DEF4C014E024DCF;
defparam prom_inst_0.INIT_RAM_15 = 256'h4E034DCD4C014E034DAD4C014E034D8D4C014E034D6D4C014E034D4D4C014E03;
defparam prom_inst_0.INIT_RAM_16 = 256'h4C014E034DCC4C014E034DAC4C014E034D8C4C014E034D6C4C014E034D4C4C01;
defparam prom_inst_0.INIT_RAM_17 = 256'h4D8A4C014E034DAB4C014E034D8B4C014E034D6B4C014E034D4B4C014E034DCB;
defparam prom_inst_0.INIT_RAM_18 = 256'h4E044D8A4C014E044DC94C014E044DCA4C014E044DCA4C014E044DAA4C014E04;
defparam prom_inst_0.INIT_RAM_19 = 256'h4C014E054DEB4C014E054D0A4C024E054D0B4C024E044DA94C014E044D894C01;
defparam prom_inst_0.INIT_RAM_1A = 256'h4D8A4C024E054D4A4C024E054D2A4C024E054D294C024E054D094C024E054DEA;
defparam prom_inst_0.INIT_RAM_1B = 256'h4E064D484C024E064DA94C024E064D894C024E064D694C024E064D494C024E06;
defparam prom_inst_0.INIT_RAM_1C = 256'h4C034E074DE94C024E074DC94C024E074DCA4C024E064D694C024E064D684C02;
defparam prom_inst_0.INIT_RAM_1D = 256'h4DE74C024E074DC74C024E074DA74C024E074DE84C024E074DC84C024E074D09;
defparam prom_inst_0.INIT_RAM_1E = 256'h61DB5D8B5C745B005808560E54C75338524751A850804F014E074D074C034E07;
defparam prom_inst_0.INIT_RAM_1F = 256'h7160700D73F06F186E506D8B6CAF6BB06AA8690068B067A8650464C0638662B8;

endmodule //Gowin_pROM
