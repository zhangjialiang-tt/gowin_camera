//Copyright (C)2014-2025 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.11.03 (64-bit)
//Part Number: GW2ANR-LV18QN88C8/I7
//Device: GW2ANR-18
//Device Version: C
//Created Time: Fri Nov  7 17:27:44 2025

module usb_retrans_ram (dout, wre, wad, di, rad, clk);

output [7:0] dout;
input wre;
input [8:0] wad;
input [7:0] di;
input [8:0] rad;
input clk;

wire wad4_inv;
wire wad5_inv;
wire wad6_inv;
wire lut_f_0;
wire wad7_inv;
wire wad8_inv;
wire lut_f_1;
wire lut_f_2;
wire lut_f_3;
wire lut_f_4;
wire lut_f_5;
wire lut_f_6;
wire lut_f_7;
wire lut_f_8;
wire lut_f_9;
wire lut_f_10;
wire lut_f_11;
wire lut_f_12;
wire lut_f_13;
wire lut_f_14;
wire lut_f_15;
wire lut_f_16;
wire lut_f_17;
wire lut_f_18;
wire lut_f_19;
wire lut_f_20;
wire lut_f_21;
wire lut_f_22;
wire lut_f_23;
wire lut_f_24;
wire lut_f_25;
wire lut_f_26;
wire lut_f_27;
wire lut_f_28;
wire lut_f_29;
wire lut_f_30;
wire lut_f_31;
wire lut_f_32;
wire lut_f_33;
wire lut_f_34;
wire lut_f_35;
wire lut_f_36;
wire lut_f_37;
wire lut_f_38;
wire lut_f_39;
wire lut_f_40;
wire lut_f_41;
wire lut_f_42;
wire lut_f_43;
wire lut_f_44;
wire lut_f_45;
wire lut_f_46;
wire lut_f_47;
wire lut_f_48;
wire lut_f_49;
wire lut_f_50;
wire lut_f_51;
wire lut_f_52;
wire lut_f_53;
wire lut_f_54;
wire lut_f_55;
wire lut_f_56;
wire lut_f_57;
wire lut_f_58;
wire lut_f_59;
wire lut_f_60;
wire lut_f_61;
wire lut_f_62;
wire lut_f_63;
wire [3:0] ram16sdp_inst_0_dout;
wire [7:4] ram16sdp_inst_1_dout;
wire [3:0] ram16sdp_inst_2_dout;
wire [7:4] ram16sdp_inst_3_dout;
wire [3:0] ram16sdp_inst_4_dout;
wire [7:4] ram16sdp_inst_5_dout;
wire [3:0] ram16sdp_inst_6_dout;
wire [7:4] ram16sdp_inst_7_dout;
wire [3:0] ram16sdp_inst_8_dout;
wire [7:4] ram16sdp_inst_9_dout;
wire [3:0] ram16sdp_inst_10_dout;
wire [7:4] ram16sdp_inst_11_dout;
wire [3:0] ram16sdp_inst_12_dout;
wire [7:4] ram16sdp_inst_13_dout;
wire [3:0] ram16sdp_inst_14_dout;
wire [7:4] ram16sdp_inst_15_dout;
wire [3:0] ram16sdp_inst_16_dout;
wire [7:4] ram16sdp_inst_17_dout;
wire [3:0] ram16sdp_inst_18_dout;
wire [7:4] ram16sdp_inst_19_dout;
wire [3:0] ram16sdp_inst_20_dout;
wire [7:4] ram16sdp_inst_21_dout;
wire [3:0] ram16sdp_inst_22_dout;
wire [7:4] ram16sdp_inst_23_dout;
wire [3:0] ram16sdp_inst_24_dout;
wire [7:4] ram16sdp_inst_25_dout;
wire [3:0] ram16sdp_inst_26_dout;
wire [7:4] ram16sdp_inst_27_dout;
wire [3:0] ram16sdp_inst_28_dout;
wire [7:4] ram16sdp_inst_29_dout;
wire [3:0] ram16sdp_inst_30_dout;
wire [7:4] ram16sdp_inst_31_dout;
wire [3:0] ram16sdp_inst_32_dout;
wire [7:4] ram16sdp_inst_33_dout;
wire [3:0] ram16sdp_inst_34_dout;
wire [7:4] ram16sdp_inst_35_dout;
wire [3:0] ram16sdp_inst_36_dout;
wire [7:4] ram16sdp_inst_37_dout;
wire [3:0] ram16sdp_inst_38_dout;
wire [7:4] ram16sdp_inst_39_dout;
wire [3:0] ram16sdp_inst_40_dout;
wire [7:4] ram16sdp_inst_41_dout;
wire [3:0] ram16sdp_inst_42_dout;
wire [7:4] ram16sdp_inst_43_dout;
wire [3:0] ram16sdp_inst_44_dout;
wire [7:4] ram16sdp_inst_45_dout;
wire [3:0] ram16sdp_inst_46_dout;
wire [7:4] ram16sdp_inst_47_dout;
wire [3:0] ram16sdp_inst_48_dout;
wire [7:4] ram16sdp_inst_49_dout;
wire [3:0] ram16sdp_inst_50_dout;
wire [7:4] ram16sdp_inst_51_dout;
wire [3:0] ram16sdp_inst_52_dout;
wire [7:4] ram16sdp_inst_53_dout;
wire [3:0] ram16sdp_inst_54_dout;
wire [7:4] ram16sdp_inst_55_dout;
wire [3:0] ram16sdp_inst_56_dout;
wire [7:4] ram16sdp_inst_57_dout;
wire [3:0] ram16sdp_inst_58_dout;
wire [7:4] ram16sdp_inst_59_dout;
wire [3:0] ram16sdp_inst_60_dout;
wire [7:4] ram16sdp_inst_61_dout;
wire [3:0] ram16sdp_inst_62_dout;
wire [7:4] ram16sdp_inst_63_dout;
wire mux_o_0;
wire mux_o_1;
wire mux_o_2;
wire mux_o_3;
wire mux_o_4;
wire mux_o_5;
wire mux_o_6;
wire mux_o_7;
wire mux_o_8;
wire mux_o_9;
wire mux_o_10;
wire mux_o_11;
wire mux_o_12;
wire mux_o_13;
wire mux_o_14;
wire mux_o_15;
wire mux_o_16;
wire mux_o_17;
wire mux_o_18;
wire mux_o_19;
wire mux_o_20;
wire mux_o_21;
wire mux_o_22;
wire mux_o_23;
wire mux_o_24;
wire mux_o_25;
wire mux_o_26;
wire mux_o_27;
wire mux_o_28;
wire mux_o_29;
wire mux_o_31;
wire mux_o_32;
wire mux_o_33;
wire mux_o_34;
wire mux_o_35;
wire mux_o_36;
wire mux_o_37;
wire mux_o_38;
wire mux_o_39;
wire mux_o_40;
wire mux_o_41;
wire mux_o_42;
wire mux_o_43;
wire mux_o_44;
wire mux_o_45;
wire mux_o_46;
wire mux_o_47;
wire mux_o_48;
wire mux_o_49;
wire mux_o_50;
wire mux_o_51;
wire mux_o_52;
wire mux_o_53;
wire mux_o_54;
wire mux_o_55;
wire mux_o_56;
wire mux_o_57;
wire mux_o_58;
wire mux_o_59;
wire mux_o_60;
wire mux_o_62;
wire mux_o_63;
wire mux_o_64;
wire mux_o_65;
wire mux_o_66;
wire mux_o_67;
wire mux_o_68;
wire mux_o_69;
wire mux_o_70;
wire mux_o_71;
wire mux_o_72;
wire mux_o_73;
wire mux_o_74;
wire mux_o_75;
wire mux_o_76;
wire mux_o_77;
wire mux_o_78;
wire mux_o_79;
wire mux_o_80;
wire mux_o_81;
wire mux_o_82;
wire mux_o_83;
wire mux_o_84;
wire mux_o_85;
wire mux_o_86;
wire mux_o_87;
wire mux_o_88;
wire mux_o_89;
wire mux_o_90;
wire mux_o_91;
wire mux_o_93;
wire mux_o_94;
wire mux_o_95;
wire mux_o_96;
wire mux_o_97;
wire mux_o_98;
wire mux_o_99;
wire mux_o_100;
wire mux_o_101;
wire mux_o_102;
wire mux_o_103;
wire mux_o_104;
wire mux_o_105;
wire mux_o_106;
wire mux_o_107;
wire mux_o_108;
wire mux_o_109;
wire mux_o_110;
wire mux_o_111;
wire mux_o_112;
wire mux_o_113;
wire mux_o_114;
wire mux_o_115;
wire mux_o_116;
wire mux_o_117;
wire mux_o_118;
wire mux_o_119;
wire mux_o_120;
wire mux_o_121;
wire mux_o_122;
wire mux_o_124;
wire mux_o_125;
wire mux_o_126;
wire mux_o_127;
wire mux_o_128;
wire mux_o_129;
wire mux_o_130;
wire mux_o_131;
wire mux_o_132;
wire mux_o_133;
wire mux_o_134;
wire mux_o_135;
wire mux_o_136;
wire mux_o_137;
wire mux_o_138;
wire mux_o_139;
wire mux_o_140;
wire mux_o_141;
wire mux_o_142;
wire mux_o_143;
wire mux_o_144;
wire mux_o_145;
wire mux_o_146;
wire mux_o_147;
wire mux_o_148;
wire mux_o_149;
wire mux_o_150;
wire mux_o_151;
wire mux_o_152;
wire mux_o_153;
wire mux_o_155;
wire mux_o_156;
wire mux_o_157;
wire mux_o_158;
wire mux_o_159;
wire mux_o_160;
wire mux_o_161;
wire mux_o_162;
wire mux_o_163;
wire mux_o_164;
wire mux_o_165;
wire mux_o_166;
wire mux_o_167;
wire mux_o_168;
wire mux_o_169;
wire mux_o_170;
wire mux_o_171;
wire mux_o_172;
wire mux_o_173;
wire mux_o_174;
wire mux_o_175;
wire mux_o_176;
wire mux_o_177;
wire mux_o_178;
wire mux_o_179;
wire mux_o_180;
wire mux_o_181;
wire mux_o_182;
wire mux_o_183;
wire mux_o_184;
wire mux_o_186;
wire mux_o_187;
wire mux_o_188;
wire mux_o_189;
wire mux_o_190;
wire mux_o_191;
wire mux_o_192;
wire mux_o_193;
wire mux_o_194;
wire mux_o_195;
wire mux_o_196;
wire mux_o_197;
wire mux_o_198;
wire mux_o_199;
wire mux_o_200;
wire mux_o_201;
wire mux_o_202;
wire mux_o_203;
wire mux_o_204;
wire mux_o_205;
wire mux_o_206;
wire mux_o_207;
wire mux_o_208;
wire mux_o_209;
wire mux_o_210;
wire mux_o_211;
wire mux_o_212;
wire mux_o_213;
wire mux_o_214;
wire mux_o_215;
wire mux_o_217;
wire mux_o_218;
wire mux_o_219;
wire mux_o_220;
wire mux_o_221;
wire mux_o_222;
wire mux_o_223;
wire mux_o_224;
wire mux_o_225;
wire mux_o_226;
wire mux_o_227;
wire mux_o_228;
wire mux_o_229;
wire mux_o_230;
wire mux_o_231;
wire mux_o_232;
wire mux_o_233;
wire mux_o_234;
wire mux_o_235;
wire mux_o_236;
wire mux_o_237;
wire mux_o_238;
wire mux_o_239;
wire mux_o_240;
wire mux_o_241;
wire mux_o_242;
wire mux_o_243;
wire mux_o_244;
wire mux_o_245;
wire mux_o_246;
wire gw_vcc;

assign gw_vcc = 1'b1;

INV inv_inst_0 (.I(wad[4]), .O(wad4_inv));

INV inv_inst_1 (.I(wad[5]), .O(wad5_inv));

INV inv_inst_2 (.I(wad[6]), .O(wad6_inv));

INV inv_inst_3 (.I(wad[7]), .O(wad7_inv));

INV inv_inst_4 (.I(wad[8]), .O(wad8_inv));

LUT4 lut_inst_0 (
  .F(lut_f_0),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_0.INIT = 16'h8000;
LUT4 lut_inst_1 (
  .F(lut_f_1),
  .I0(lut_f_0),
  .I1(wad7_inv),
  .I2(wad8_inv),
  .I3(gw_vcc)
);
defparam lut_inst_1.INIT = 16'h8000;
LUT4 lut_inst_2 (
  .F(lut_f_2),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_2.INIT = 16'h8000;
LUT4 lut_inst_3 (
  .F(lut_f_3),
  .I0(lut_f_2),
  .I1(wad7_inv),
  .I2(wad8_inv),
  .I3(gw_vcc)
);
defparam lut_inst_3.INIT = 16'h8000;
LUT4 lut_inst_4 (
  .F(lut_f_4),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_4.INIT = 16'h8000;
LUT4 lut_inst_5 (
  .F(lut_f_5),
  .I0(lut_f_4),
  .I1(wad7_inv),
  .I2(wad8_inv),
  .I3(gw_vcc)
);
defparam lut_inst_5.INIT = 16'h8000;
LUT4 lut_inst_6 (
  .F(lut_f_6),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_6.INIT = 16'h8000;
LUT4 lut_inst_7 (
  .F(lut_f_7),
  .I0(lut_f_6),
  .I1(wad7_inv),
  .I2(wad8_inv),
  .I3(gw_vcc)
);
defparam lut_inst_7.INIT = 16'h8000;
LUT4 lut_inst_8 (
  .F(lut_f_8),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_8.INIT = 16'h8000;
LUT4 lut_inst_9 (
  .F(lut_f_9),
  .I0(lut_f_8),
  .I1(wad7_inv),
  .I2(wad8_inv),
  .I3(gw_vcc)
);
defparam lut_inst_9.INIT = 16'h8000;
LUT4 lut_inst_10 (
  .F(lut_f_10),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_10.INIT = 16'h8000;
LUT4 lut_inst_11 (
  .F(lut_f_11),
  .I0(lut_f_10),
  .I1(wad7_inv),
  .I2(wad8_inv),
  .I3(gw_vcc)
);
defparam lut_inst_11.INIT = 16'h8000;
LUT4 lut_inst_12 (
  .F(lut_f_12),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_12.INIT = 16'h8000;
LUT4 lut_inst_13 (
  .F(lut_f_13),
  .I0(lut_f_12),
  .I1(wad7_inv),
  .I2(wad8_inv),
  .I3(gw_vcc)
);
defparam lut_inst_13.INIT = 16'h8000;
LUT4 lut_inst_14 (
  .F(lut_f_14),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_14.INIT = 16'h8000;
LUT4 lut_inst_15 (
  .F(lut_f_15),
  .I0(lut_f_14),
  .I1(wad7_inv),
  .I2(wad8_inv),
  .I3(gw_vcc)
);
defparam lut_inst_15.INIT = 16'h8000;
LUT4 lut_inst_16 (
  .F(lut_f_16),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_16.INIT = 16'h8000;
LUT4 lut_inst_17 (
  .F(lut_f_17),
  .I0(lut_f_16),
  .I1(wad[7]),
  .I2(wad8_inv),
  .I3(gw_vcc)
);
defparam lut_inst_17.INIT = 16'h8000;
LUT4 lut_inst_18 (
  .F(lut_f_18),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_18.INIT = 16'h8000;
LUT4 lut_inst_19 (
  .F(lut_f_19),
  .I0(lut_f_18),
  .I1(wad[7]),
  .I2(wad8_inv),
  .I3(gw_vcc)
);
defparam lut_inst_19.INIT = 16'h8000;
LUT4 lut_inst_20 (
  .F(lut_f_20),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_20.INIT = 16'h8000;
LUT4 lut_inst_21 (
  .F(lut_f_21),
  .I0(lut_f_20),
  .I1(wad[7]),
  .I2(wad8_inv),
  .I3(gw_vcc)
);
defparam lut_inst_21.INIT = 16'h8000;
LUT4 lut_inst_22 (
  .F(lut_f_22),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_22.INIT = 16'h8000;
LUT4 lut_inst_23 (
  .F(lut_f_23),
  .I0(lut_f_22),
  .I1(wad[7]),
  .I2(wad8_inv),
  .I3(gw_vcc)
);
defparam lut_inst_23.INIT = 16'h8000;
LUT4 lut_inst_24 (
  .F(lut_f_24),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_24.INIT = 16'h8000;
LUT4 lut_inst_25 (
  .F(lut_f_25),
  .I0(lut_f_24),
  .I1(wad[7]),
  .I2(wad8_inv),
  .I3(gw_vcc)
);
defparam lut_inst_25.INIT = 16'h8000;
LUT4 lut_inst_26 (
  .F(lut_f_26),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_26.INIT = 16'h8000;
LUT4 lut_inst_27 (
  .F(lut_f_27),
  .I0(lut_f_26),
  .I1(wad[7]),
  .I2(wad8_inv),
  .I3(gw_vcc)
);
defparam lut_inst_27.INIT = 16'h8000;
LUT4 lut_inst_28 (
  .F(lut_f_28),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_28.INIT = 16'h8000;
LUT4 lut_inst_29 (
  .F(lut_f_29),
  .I0(lut_f_28),
  .I1(wad[7]),
  .I2(wad8_inv),
  .I3(gw_vcc)
);
defparam lut_inst_29.INIT = 16'h8000;
LUT4 lut_inst_30 (
  .F(lut_f_30),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_30.INIT = 16'h8000;
LUT4 lut_inst_31 (
  .F(lut_f_31),
  .I0(lut_f_30),
  .I1(wad[7]),
  .I2(wad8_inv),
  .I3(gw_vcc)
);
defparam lut_inst_31.INIT = 16'h8000;
LUT4 lut_inst_32 (
  .F(lut_f_32),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_32.INIT = 16'h8000;
LUT4 lut_inst_33 (
  .F(lut_f_33),
  .I0(lut_f_32),
  .I1(wad7_inv),
  .I2(wad[8]),
  .I3(gw_vcc)
);
defparam lut_inst_33.INIT = 16'h8000;
LUT4 lut_inst_34 (
  .F(lut_f_34),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_34.INIT = 16'h8000;
LUT4 lut_inst_35 (
  .F(lut_f_35),
  .I0(lut_f_34),
  .I1(wad7_inv),
  .I2(wad[8]),
  .I3(gw_vcc)
);
defparam lut_inst_35.INIT = 16'h8000;
LUT4 lut_inst_36 (
  .F(lut_f_36),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_36.INIT = 16'h8000;
LUT4 lut_inst_37 (
  .F(lut_f_37),
  .I0(lut_f_36),
  .I1(wad7_inv),
  .I2(wad[8]),
  .I3(gw_vcc)
);
defparam lut_inst_37.INIT = 16'h8000;
LUT4 lut_inst_38 (
  .F(lut_f_38),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_38.INIT = 16'h8000;
LUT4 lut_inst_39 (
  .F(lut_f_39),
  .I0(lut_f_38),
  .I1(wad7_inv),
  .I2(wad[8]),
  .I3(gw_vcc)
);
defparam lut_inst_39.INIT = 16'h8000;
LUT4 lut_inst_40 (
  .F(lut_f_40),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_40.INIT = 16'h8000;
LUT4 lut_inst_41 (
  .F(lut_f_41),
  .I0(lut_f_40),
  .I1(wad7_inv),
  .I2(wad[8]),
  .I3(gw_vcc)
);
defparam lut_inst_41.INIT = 16'h8000;
LUT4 lut_inst_42 (
  .F(lut_f_42),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_42.INIT = 16'h8000;
LUT4 lut_inst_43 (
  .F(lut_f_43),
  .I0(lut_f_42),
  .I1(wad7_inv),
  .I2(wad[8]),
  .I3(gw_vcc)
);
defparam lut_inst_43.INIT = 16'h8000;
LUT4 lut_inst_44 (
  .F(lut_f_44),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_44.INIT = 16'h8000;
LUT4 lut_inst_45 (
  .F(lut_f_45),
  .I0(lut_f_44),
  .I1(wad7_inv),
  .I2(wad[8]),
  .I3(gw_vcc)
);
defparam lut_inst_45.INIT = 16'h8000;
LUT4 lut_inst_46 (
  .F(lut_f_46),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_46.INIT = 16'h8000;
LUT4 lut_inst_47 (
  .F(lut_f_47),
  .I0(lut_f_46),
  .I1(wad7_inv),
  .I2(wad[8]),
  .I3(gw_vcc)
);
defparam lut_inst_47.INIT = 16'h8000;
LUT4 lut_inst_48 (
  .F(lut_f_48),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_48.INIT = 16'h8000;
LUT4 lut_inst_49 (
  .F(lut_f_49),
  .I0(lut_f_48),
  .I1(wad[7]),
  .I2(wad[8]),
  .I3(gw_vcc)
);
defparam lut_inst_49.INIT = 16'h8000;
LUT4 lut_inst_50 (
  .F(lut_f_50),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_50.INIT = 16'h8000;
LUT4 lut_inst_51 (
  .F(lut_f_51),
  .I0(lut_f_50),
  .I1(wad[7]),
  .I2(wad[8]),
  .I3(gw_vcc)
);
defparam lut_inst_51.INIT = 16'h8000;
LUT4 lut_inst_52 (
  .F(lut_f_52),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_52.INIT = 16'h8000;
LUT4 lut_inst_53 (
  .F(lut_f_53),
  .I0(lut_f_52),
  .I1(wad[7]),
  .I2(wad[8]),
  .I3(gw_vcc)
);
defparam lut_inst_53.INIT = 16'h8000;
LUT4 lut_inst_54 (
  .F(lut_f_54),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_54.INIT = 16'h8000;
LUT4 lut_inst_55 (
  .F(lut_f_55),
  .I0(lut_f_54),
  .I1(wad[7]),
  .I2(wad[8]),
  .I3(gw_vcc)
);
defparam lut_inst_55.INIT = 16'h8000;
LUT4 lut_inst_56 (
  .F(lut_f_56),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_56.INIT = 16'h8000;
LUT4 lut_inst_57 (
  .F(lut_f_57),
  .I0(lut_f_56),
  .I1(wad[7]),
  .I2(wad[8]),
  .I3(gw_vcc)
);
defparam lut_inst_57.INIT = 16'h8000;
LUT4 lut_inst_58 (
  .F(lut_f_58),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_58.INIT = 16'h8000;
LUT4 lut_inst_59 (
  .F(lut_f_59),
  .I0(lut_f_58),
  .I1(wad[7]),
  .I2(wad[8]),
  .I3(gw_vcc)
);
defparam lut_inst_59.INIT = 16'h8000;
LUT4 lut_inst_60 (
  .F(lut_f_60),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_60.INIT = 16'h8000;
LUT4 lut_inst_61 (
  .F(lut_f_61),
  .I0(lut_f_60),
  .I1(wad[7]),
  .I2(wad[8]),
  .I3(gw_vcc)
);
defparam lut_inst_61.INIT = 16'h8000;
LUT4 lut_inst_62 (
  .F(lut_f_62),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_62.INIT = 16'h8000;
LUT4 lut_inst_63 (
  .F(lut_f_63),
  .I0(lut_f_62),
  .I1(wad[7]),
  .I2(wad[8]),
  .I3(gw_vcc)
);
defparam lut_inst_63.INIT = 16'h8000;
RAM16SDP4 ram16sdp_inst_0 (
    .DO(ram16sdp_inst_0_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16sdp_inst_0.INIT_0 = 16'h0000;
defparam ram16sdp_inst_0.INIT_1 = 16'h0000;
defparam ram16sdp_inst_0.INIT_2 = 16'h0000;
defparam ram16sdp_inst_0.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_1 (
    .DO(ram16sdp_inst_1_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16sdp_inst_1.INIT_0 = 16'h0000;
defparam ram16sdp_inst_1.INIT_1 = 16'h0000;
defparam ram16sdp_inst_1.INIT_2 = 16'h0000;
defparam ram16sdp_inst_1.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_2 (
    .DO(ram16sdp_inst_2_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_3),
    .CLK(clk)
);

defparam ram16sdp_inst_2.INIT_0 = 16'h0000;
defparam ram16sdp_inst_2.INIT_1 = 16'h0000;
defparam ram16sdp_inst_2.INIT_2 = 16'h0000;
defparam ram16sdp_inst_2.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_3 (
    .DO(ram16sdp_inst_3_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_3),
    .CLK(clk)
);

defparam ram16sdp_inst_3.INIT_0 = 16'h0000;
defparam ram16sdp_inst_3.INIT_1 = 16'h0000;
defparam ram16sdp_inst_3.INIT_2 = 16'h0000;
defparam ram16sdp_inst_3.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_4 (
    .DO(ram16sdp_inst_4_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_5),
    .CLK(clk)
);

defparam ram16sdp_inst_4.INIT_0 = 16'h0000;
defparam ram16sdp_inst_4.INIT_1 = 16'h0000;
defparam ram16sdp_inst_4.INIT_2 = 16'h0000;
defparam ram16sdp_inst_4.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_5 (
    .DO(ram16sdp_inst_5_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_5),
    .CLK(clk)
);

defparam ram16sdp_inst_5.INIT_0 = 16'h0000;
defparam ram16sdp_inst_5.INIT_1 = 16'h0000;
defparam ram16sdp_inst_5.INIT_2 = 16'h0000;
defparam ram16sdp_inst_5.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_6 (
    .DO(ram16sdp_inst_6_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_7),
    .CLK(clk)
);

defparam ram16sdp_inst_6.INIT_0 = 16'h0000;
defparam ram16sdp_inst_6.INIT_1 = 16'h0000;
defparam ram16sdp_inst_6.INIT_2 = 16'h0000;
defparam ram16sdp_inst_6.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_7 (
    .DO(ram16sdp_inst_7_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_7),
    .CLK(clk)
);

defparam ram16sdp_inst_7.INIT_0 = 16'h0000;
defparam ram16sdp_inst_7.INIT_1 = 16'h0000;
defparam ram16sdp_inst_7.INIT_2 = 16'h0000;
defparam ram16sdp_inst_7.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_8 (
    .DO(ram16sdp_inst_8_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_9),
    .CLK(clk)
);

defparam ram16sdp_inst_8.INIT_0 = 16'h0000;
defparam ram16sdp_inst_8.INIT_1 = 16'h0000;
defparam ram16sdp_inst_8.INIT_2 = 16'h0000;
defparam ram16sdp_inst_8.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_9 (
    .DO(ram16sdp_inst_9_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_9),
    .CLK(clk)
);

defparam ram16sdp_inst_9.INIT_0 = 16'h0000;
defparam ram16sdp_inst_9.INIT_1 = 16'h0000;
defparam ram16sdp_inst_9.INIT_2 = 16'h0000;
defparam ram16sdp_inst_9.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_10 (
    .DO(ram16sdp_inst_10_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_11),
    .CLK(clk)
);

defparam ram16sdp_inst_10.INIT_0 = 16'h0000;
defparam ram16sdp_inst_10.INIT_1 = 16'h0000;
defparam ram16sdp_inst_10.INIT_2 = 16'h0000;
defparam ram16sdp_inst_10.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_11 (
    .DO(ram16sdp_inst_11_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_11),
    .CLK(clk)
);

defparam ram16sdp_inst_11.INIT_0 = 16'h0000;
defparam ram16sdp_inst_11.INIT_1 = 16'h0000;
defparam ram16sdp_inst_11.INIT_2 = 16'h0000;
defparam ram16sdp_inst_11.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_12 (
    .DO(ram16sdp_inst_12_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_13),
    .CLK(clk)
);

defparam ram16sdp_inst_12.INIT_0 = 16'h0000;
defparam ram16sdp_inst_12.INIT_1 = 16'h0000;
defparam ram16sdp_inst_12.INIT_2 = 16'h0000;
defparam ram16sdp_inst_12.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_13 (
    .DO(ram16sdp_inst_13_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_13),
    .CLK(clk)
);

defparam ram16sdp_inst_13.INIT_0 = 16'h0000;
defparam ram16sdp_inst_13.INIT_1 = 16'h0000;
defparam ram16sdp_inst_13.INIT_2 = 16'h0000;
defparam ram16sdp_inst_13.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_14 (
    .DO(ram16sdp_inst_14_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_15),
    .CLK(clk)
);

defparam ram16sdp_inst_14.INIT_0 = 16'h0000;
defparam ram16sdp_inst_14.INIT_1 = 16'h0000;
defparam ram16sdp_inst_14.INIT_2 = 16'h0000;
defparam ram16sdp_inst_14.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_15 (
    .DO(ram16sdp_inst_15_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_15),
    .CLK(clk)
);

defparam ram16sdp_inst_15.INIT_0 = 16'h0000;
defparam ram16sdp_inst_15.INIT_1 = 16'h0000;
defparam ram16sdp_inst_15.INIT_2 = 16'h0000;
defparam ram16sdp_inst_15.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_16 (
    .DO(ram16sdp_inst_16_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_17),
    .CLK(clk)
);

defparam ram16sdp_inst_16.INIT_0 = 16'h0000;
defparam ram16sdp_inst_16.INIT_1 = 16'h0000;
defparam ram16sdp_inst_16.INIT_2 = 16'h0000;
defparam ram16sdp_inst_16.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_17 (
    .DO(ram16sdp_inst_17_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_17),
    .CLK(clk)
);

defparam ram16sdp_inst_17.INIT_0 = 16'h0000;
defparam ram16sdp_inst_17.INIT_1 = 16'h0000;
defparam ram16sdp_inst_17.INIT_2 = 16'h0000;
defparam ram16sdp_inst_17.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_18 (
    .DO(ram16sdp_inst_18_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_19),
    .CLK(clk)
);

defparam ram16sdp_inst_18.INIT_0 = 16'h0000;
defparam ram16sdp_inst_18.INIT_1 = 16'h0000;
defparam ram16sdp_inst_18.INIT_2 = 16'h0000;
defparam ram16sdp_inst_18.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_19 (
    .DO(ram16sdp_inst_19_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_19),
    .CLK(clk)
);

defparam ram16sdp_inst_19.INIT_0 = 16'h0000;
defparam ram16sdp_inst_19.INIT_1 = 16'h0000;
defparam ram16sdp_inst_19.INIT_2 = 16'h0000;
defparam ram16sdp_inst_19.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_20 (
    .DO(ram16sdp_inst_20_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_21),
    .CLK(clk)
);

defparam ram16sdp_inst_20.INIT_0 = 16'h0000;
defparam ram16sdp_inst_20.INIT_1 = 16'h0000;
defparam ram16sdp_inst_20.INIT_2 = 16'h0000;
defparam ram16sdp_inst_20.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_21 (
    .DO(ram16sdp_inst_21_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_21),
    .CLK(clk)
);

defparam ram16sdp_inst_21.INIT_0 = 16'h0000;
defparam ram16sdp_inst_21.INIT_1 = 16'h0000;
defparam ram16sdp_inst_21.INIT_2 = 16'h0000;
defparam ram16sdp_inst_21.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_22 (
    .DO(ram16sdp_inst_22_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_23),
    .CLK(clk)
);

defparam ram16sdp_inst_22.INIT_0 = 16'h0000;
defparam ram16sdp_inst_22.INIT_1 = 16'h0000;
defparam ram16sdp_inst_22.INIT_2 = 16'h0000;
defparam ram16sdp_inst_22.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_23 (
    .DO(ram16sdp_inst_23_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_23),
    .CLK(clk)
);

defparam ram16sdp_inst_23.INIT_0 = 16'h0000;
defparam ram16sdp_inst_23.INIT_1 = 16'h0000;
defparam ram16sdp_inst_23.INIT_2 = 16'h0000;
defparam ram16sdp_inst_23.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_24 (
    .DO(ram16sdp_inst_24_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_25),
    .CLK(clk)
);

defparam ram16sdp_inst_24.INIT_0 = 16'h0000;
defparam ram16sdp_inst_24.INIT_1 = 16'h0000;
defparam ram16sdp_inst_24.INIT_2 = 16'h0000;
defparam ram16sdp_inst_24.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_25 (
    .DO(ram16sdp_inst_25_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_25),
    .CLK(clk)
);

defparam ram16sdp_inst_25.INIT_0 = 16'h0000;
defparam ram16sdp_inst_25.INIT_1 = 16'h0000;
defparam ram16sdp_inst_25.INIT_2 = 16'h0000;
defparam ram16sdp_inst_25.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_26 (
    .DO(ram16sdp_inst_26_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_27),
    .CLK(clk)
);

defparam ram16sdp_inst_26.INIT_0 = 16'h0000;
defparam ram16sdp_inst_26.INIT_1 = 16'h0000;
defparam ram16sdp_inst_26.INIT_2 = 16'h0000;
defparam ram16sdp_inst_26.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_27 (
    .DO(ram16sdp_inst_27_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_27),
    .CLK(clk)
);

defparam ram16sdp_inst_27.INIT_0 = 16'h0000;
defparam ram16sdp_inst_27.INIT_1 = 16'h0000;
defparam ram16sdp_inst_27.INIT_2 = 16'h0000;
defparam ram16sdp_inst_27.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_28 (
    .DO(ram16sdp_inst_28_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_29),
    .CLK(clk)
);

defparam ram16sdp_inst_28.INIT_0 = 16'h0000;
defparam ram16sdp_inst_28.INIT_1 = 16'h0000;
defparam ram16sdp_inst_28.INIT_2 = 16'h0000;
defparam ram16sdp_inst_28.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_29 (
    .DO(ram16sdp_inst_29_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_29),
    .CLK(clk)
);

defparam ram16sdp_inst_29.INIT_0 = 16'h0000;
defparam ram16sdp_inst_29.INIT_1 = 16'h0000;
defparam ram16sdp_inst_29.INIT_2 = 16'h0000;
defparam ram16sdp_inst_29.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_30 (
    .DO(ram16sdp_inst_30_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_31),
    .CLK(clk)
);

defparam ram16sdp_inst_30.INIT_0 = 16'h0000;
defparam ram16sdp_inst_30.INIT_1 = 16'h0000;
defparam ram16sdp_inst_30.INIT_2 = 16'h0000;
defparam ram16sdp_inst_30.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_31 (
    .DO(ram16sdp_inst_31_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_31),
    .CLK(clk)
);

defparam ram16sdp_inst_31.INIT_0 = 16'h0000;
defparam ram16sdp_inst_31.INIT_1 = 16'h0000;
defparam ram16sdp_inst_31.INIT_2 = 16'h0000;
defparam ram16sdp_inst_31.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_32 (
    .DO(ram16sdp_inst_32_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_33),
    .CLK(clk)
);

defparam ram16sdp_inst_32.INIT_0 = 16'h0000;
defparam ram16sdp_inst_32.INIT_1 = 16'h0000;
defparam ram16sdp_inst_32.INIT_2 = 16'h0000;
defparam ram16sdp_inst_32.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_33 (
    .DO(ram16sdp_inst_33_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_33),
    .CLK(clk)
);

defparam ram16sdp_inst_33.INIT_0 = 16'h0000;
defparam ram16sdp_inst_33.INIT_1 = 16'h0000;
defparam ram16sdp_inst_33.INIT_2 = 16'h0000;
defparam ram16sdp_inst_33.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_34 (
    .DO(ram16sdp_inst_34_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_35),
    .CLK(clk)
);

defparam ram16sdp_inst_34.INIT_0 = 16'h0000;
defparam ram16sdp_inst_34.INIT_1 = 16'h0000;
defparam ram16sdp_inst_34.INIT_2 = 16'h0000;
defparam ram16sdp_inst_34.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_35 (
    .DO(ram16sdp_inst_35_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_35),
    .CLK(clk)
);

defparam ram16sdp_inst_35.INIT_0 = 16'h0000;
defparam ram16sdp_inst_35.INIT_1 = 16'h0000;
defparam ram16sdp_inst_35.INIT_2 = 16'h0000;
defparam ram16sdp_inst_35.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_36 (
    .DO(ram16sdp_inst_36_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_37),
    .CLK(clk)
);

defparam ram16sdp_inst_36.INIT_0 = 16'h0000;
defparam ram16sdp_inst_36.INIT_1 = 16'h0000;
defparam ram16sdp_inst_36.INIT_2 = 16'h0000;
defparam ram16sdp_inst_36.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_37 (
    .DO(ram16sdp_inst_37_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_37),
    .CLK(clk)
);

defparam ram16sdp_inst_37.INIT_0 = 16'h0000;
defparam ram16sdp_inst_37.INIT_1 = 16'h0000;
defparam ram16sdp_inst_37.INIT_2 = 16'h0000;
defparam ram16sdp_inst_37.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_38 (
    .DO(ram16sdp_inst_38_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_39),
    .CLK(clk)
);

defparam ram16sdp_inst_38.INIT_0 = 16'h0000;
defparam ram16sdp_inst_38.INIT_1 = 16'h0000;
defparam ram16sdp_inst_38.INIT_2 = 16'h0000;
defparam ram16sdp_inst_38.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_39 (
    .DO(ram16sdp_inst_39_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_39),
    .CLK(clk)
);

defparam ram16sdp_inst_39.INIT_0 = 16'h0000;
defparam ram16sdp_inst_39.INIT_1 = 16'h0000;
defparam ram16sdp_inst_39.INIT_2 = 16'h0000;
defparam ram16sdp_inst_39.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_40 (
    .DO(ram16sdp_inst_40_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_41),
    .CLK(clk)
);

defparam ram16sdp_inst_40.INIT_0 = 16'h0000;
defparam ram16sdp_inst_40.INIT_1 = 16'h0000;
defparam ram16sdp_inst_40.INIT_2 = 16'h0000;
defparam ram16sdp_inst_40.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_41 (
    .DO(ram16sdp_inst_41_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_41),
    .CLK(clk)
);

defparam ram16sdp_inst_41.INIT_0 = 16'h0000;
defparam ram16sdp_inst_41.INIT_1 = 16'h0000;
defparam ram16sdp_inst_41.INIT_2 = 16'h0000;
defparam ram16sdp_inst_41.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_42 (
    .DO(ram16sdp_inst_42_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_43),
    .CLK(clk)
);

defparam ram16sdp_inst_42.INIT_0 = 16'h0000;
defparam ram16sdp_inst_42.INIT_1 = 16'h0000;
defparam ram16sdp_inst_42.INIT_2 = 16'h0000;
defparam ram16sdp_inst_42.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_43 (
    .DO(ram16sdp_inst_43_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_43),
    .CLK(clk)
);

defparam ram16sdp_inst_43.INIT_0 = 16'h0000;
defparam ram16sdp_inst_43.INIT_1 = 16'h0000;
defparam ram16sdp_inst_43.INIT_2 = 16'h0000;
defparam ram16sdp_inst_43.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_44 (
    .DO(ram16sdp_inst_44_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_45),
    .CLK(clk)
);

defparam ram16sdp_inst_44.INIT_0 = 16'h0000;
defparam ram16sdp_inst_44.INIT_1 = 16'h0000;
defparam ram16sdp_inst_44.INIT_2 = 16'h0000;
defparam ram16sdp_inst_44.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_45 (
    .DO(ram16sdp_inst_45_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_45),
    .CLK(clk)
);

defparam ram16sdp_inst_45.INIT_0 = 16'h0000;
defparam ram16sdp_inst_45.INIT_1 = 16'h0000;
defparam ram16sdp_inst_45.INIT_2 = 16'h0000;
defparam ram16sdp_inst_45.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_46 (
    .DO(ram16sdp_inst_46_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_47),
    .CLK(clk)
);

defparam ram16sdp_inst_46.INIT_0 = 16'h0000;
defparam ram16sdp_inst_46.INIT_1 = 16'h0000;
defparam ram16sdp_inst_46.INIT_2 = 16'h0000;
defparam ram16sdp_inst_46.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_47 (
    .DO(ram16sdp_inst_47_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_47),
    .CLK(clk)
);

defparam ram16sdp_inst_47.INIT_0 = 16'h0000;
defparam ram16sdp_inst_47.INIT_1 = 16'h0000;
defparam ram16sdp_inst_47.INIT_2 = 16'h0000;
defparam ram16sdp_inst_47.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_48 (
    .DO(ram16sdp_inst_48_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_49),
    .CLK(clk)
);

defparam ram16sdp_inst_48.INIT_0 = 16'h0000;
defparam ram16sdp_inst_48.INIT_1 = 16'h0000;
defparam ram16sdp_inst_48.INIT_2 = 16'h0000;
defparam ram16sdp_inst_48.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_49 (
    .DO(ram16sdp_inst_49_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_49),
    .CLK(clk)
);

defparam ram16sdp_inst_49.INIT_0 = 16'h0000;
defparam ram16sdp_inst_49.INIT_1 = 16'h0000;
defparam ram16sdp_inst_49.INIT_2 = 16'h0000;
defparam ram16sdp_inst_49.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_50 (
    .DO(ram16sdp_inst_50_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_51),
    .CLK(clk)
);

defparam ram16sdp_inst_50.INIT_0 = 16'h0000;
defparam ram16sdp_inst_50.INIT_1 = 16'h0000;
defparam ram16sdp_inst_50.INIT_2 = 16'h0000;
defparam ram16sdp_inst_50.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_51 (
    .DO(ram16sdp_inst_51_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_51),
    .CLK(clk)
);

defparam ram16sdp_inst_51.INIT_0 = 16'h0000;
defparam ram16sdp_inst_51.INIT_1 = 16'h0000;
defparam ram16sdp_inst_51.INIT_2 = 16'h0000;
defparam ram16sdp_inst_51.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_52 (
    .DO(ram16sdp_inst_52_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_53),
    .CLK(clk)
);

defparam ram16sdp_inst_52.INIT_0 = 16'h0000;
defparam ram16sdp_inst_52.INIT_1 = 16'h0000;
defparam ram16sdp_inst_52.INIT_2 = 16'h0000;
defparam ram16sdp_inst_52.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_53 (
    .DO(ram16sdp_inst_53_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_53),
    .CLK(clk)
);

defparam ram16sdp_inst_53.INIT_0 = 16'h0000;
defparam ram16sdp_inst_53.INIT_1 = 16'h0000;
defparam ram16sdp_inst_53.INIT_2 = 16'h0000;
defparam ram16sdp_inst_53.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_54 (
    .DO(ram16sdp_inst_54_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_55),
    .CLK(clk)
);

defparam ram16sdp_inst_54.INIT_0 = 16'h0000;
defparam ram16sdp_inst_54.INIT_1 = 16'h0000;
defparam ram16sdp_inst_54.INIT_2 = 16'h0000;
defparam ram16sdp_inst_54.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_55 (
    .DO(ram16sdp_inst_55_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_55),
    .CLK(clk)
);

defparam ram16sdp_inst_55.INIT_0 = 16'h0000;
defparam ram16sdp_inst_55.INIT_1 = 16'h0000;
defparam ram16sdp_inst_55.INIT_2 = 16'h0000;
defparam ram16sdp_inst_55.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_56 (
    .DO(ram16sdp_inst_56_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_57),
    .CLK(clk)
);

defparam ram16sdp_inst_56.INIT_0 = 16'h0000;
defparam ram16sdp_inst_56.INIT_1 = 16'h0000;
defparam ram16sdp_inst_56.INIT_2 = 16'h0000;
defparam ram16sdp_inst_56.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_57 (
    .DO(ram16sdp_inst_57_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_57),
    .CLK(clk)
);

defparam ram16sdp_inst_57.INIT_0 = 16'h0000;
defparam ram16sdp_inst_57.INIT_1 = 16'h0000;
defparam ram16sdp_inst_57.INIT_2 = 16'h0000;
defparam ram16sdp_inst_57.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_58 (
    .DO(ram16sdp_inst_58_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_59),
    .CLK(clk)
);

defparam ram16sdp_inst_58.INIT_0 = 16'h0000;
defparam ram16sdp_inst_58.INIT_1 = 16'h0000;
defparam ram16sdp_inst_58.INIT_2 = 16'h0000;
defparam ram16sdp_inst_58.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_59 (
    .DO(ram16sdp_inst_59_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_59),
    .CLK(clk)
);

defparam ram16sdp_inst_59.INIT_0 = 16'h0000;
defparam ram16sdp_inst_59.INIT_1 = 16'h0000;
defparam ram16sdp_inst_59.INIT_2 = 16'h0000;
defparam ram16sdp_inst_59.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_60 (
    .DO(ram16sdp_inst_60_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_61),
    .CLK(clk)
);

defparam ram16sdp_inst_60.INIT_0 = 16'h0000;
defparam ram16sdp_inst_60.INIT_1 = 16'h0000;
defparam ram16sdp_inst_60.INIT_2 = 16'h0000;
defparam ram16sdp_inst_60.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_61 (
    .DO(ram16sdp_inst_61_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_61),
    .CLK(clk)
);

defparam ram16sdp_inst_61.INIT_0 = 16'h0000;
defparam ram16sdp_inst_61.INIT_1 = 16'h0000;
defparam ram16sdp_inst_61.INIT_2 = 16'h0000;
defparam ram16sdp_inst_61.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_62 (
    .DO(ram16sdp_inst_62_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_63),
    .CLK(clk)
);

defparam ram16sdp_inst_62.INIT_0 = 16'h0000;
defparam ram16sdp_inst_62.INIT_1 = 16'h0000;
defparam ram16sdp_inst_62.INIT_2 = 16'h0000;
defparam ram16sdp_inst_62.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_63 (
    .DO(ram16sdp_inst_63_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_63),
    .CLK(clk)
);

defparam ram16sdp_inst_63.INIT_0 = 16'h0000;
defparam ram16sdp_inst_63.INIT_1 = 16'h0000;
defparam ram16sdp_inst_63.INIT_2 = 16'h0000;
defparam ram16sdp_inst_63.INIT_3 = 16'h0000;

MUX2 mux_inst_0 (
  .O(mux_o_0),
  .I0(ram16sdp_inst_0_dout[0]),
  .I1(ram16sdp_inst_2_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_1 (
  .O(mux_o_1),
  .I0(ram16sdp_inst_4_dout[0]),
  .I1(ram16sdp_inst_6_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_2 (
  .O(mux_o_2),
  .I0(ram16sdp_inst_8_dout[0]),
  .I1(ram16sdp_inst_10_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_3 (
  .O(mux_o_3),
  .I0(ram16sdp_inst_12_dout[0]),
  .I1(ram16sdp_inst_14_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_4 (
  .O(mux_o_4),
  .I0(ram16sdp_inst_16_dout[0]),
  .I1(ram16sdp_inst_18_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_5 (
  .O(mux_o_5),
  .I0(ram16sdp_inst_20_dout[0]),
  .I1(ram16sdp_inst_22_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_6 (
  .O(mux_o_6),
  .I0(ram16sdp_inst_24_dout[0]),
  .I1(ram16sdp_inst_26_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_7 (
  .O(mux_o_7),
  .I0(ram16sdp_inst_28_dout[0]),
  .I1(ram16sdp_inst_30_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_8 (
  .O(mux_o_8),
  .I0(ram16sdp_inst_32_dout[0]),
  .I1(ram16sdp_inst_34_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_9 (
  .O(mux_o_9),
  .I0(ram16sdp_inst_36_dout[0]),
  .I1(ram16sdp_inst_38_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_10 (
  .O(mux_o_10),
  .I0(ram16sdp_inst_40_dout[0]),
  .I1(ram16sdp_inst_42_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_11 (
  .O(mux_o_11),
  .I0(ram16sdp_inst_44_dout[0]),
  .I1(ram16sdp_inst_46_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_12 (
  .O(mux_o_12),
  .I0(ram16sdp_inst_48_dout[0]),
  .I1(ram16sdp_inst_50_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_13 (
  .O(mux_o_13),
  .I0(ram16sdp_inst_52_dout[0]),
  .I1(ram16sdp_inst_54_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_14 (
  .O(mux_o_14),
  .I0(ram16sdp_inst_56_dout[0]),
  .I1(ram16sdp_inst_58_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_15 (
  .O(mux_o_15),
  .I0(ram16sdp_inst_60_dout[0]),
  .I1(ram16sdp_inst_62_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_16 (
  .O(mux_o_16),
  .I0(mux_o_0),
  .I1(mux_o_1),
  .S0(rad[5])
);
MUX2 mux_inst_17 (
  .O(mux_o_17),
  .I0(mux_o_2),
  .I1(mux_o_3),
  .S0(rad[5])
);
MUX2 mux_inst_18 (
  .O(mux_o_18),
  .I0(mux_o_4),
  .I1(mux_o_5),
  .S0(rad[5])
);
MUX2 mux_inst_19 (
  .O(mux_o_19),
  .I0(mux_o_6),
  .I1(mux_o_7),
  .S0(rad[5])
);
MUX2 mux_inst_20 (
  .O(mux_o_20),
  .I0(mux_o_8),
  .I1(mux_o_9),
  .S0(rad[5])
);
MUX2 mux_inst_21 (
  .O(mux_o_21),
  .I0(mux_o_10),
  .I1(mux_o_11),
  .S0(rad[5])
);
MUX2 mux_inst_22 (
  .O(mux_o_22),
  .I0(mux_o_12),
  .I1(mux_o_13),
  .S0(rad[5])
);
MUX2 mux_inst_23 (
  .O(mux_o_23),
  .I0(mux_o_14),
  .I1(mux_o_15),
  .S0(rad[5])
);
MUX2 mux_inst_24 (
  .O(mux_o_24),
  .I0(mux_o_16),
  .I1(mux_o_17),
  .S0(rad[6])
);
MUX2 mux_inst_25 (
  .O(mux_o_25),
  .I0(mux_o_18),
  .I1(mux_o_19),
  .S0(rad[6])
);
MUX2 mux_inst_26 (
  .O(mux_o_26),
  .I0(mux_o_20),
  .I1(mux_o_21),
  .S0(rad[6])
);
MUX2 mux_inst_27 (
  .O(mux_o_27),
  .I0(mux_o_22),
  .I1(mux_o_23),
  .S0(rad[6])
);
MUX2 mux_inst_28 (
  .O(mux_o_28),
  .I0(mux_o_24),
  .I1(mux_o_25),
  .S0(rad[7])
);
MUX2 mux_inst_29 (
  .O(mux_o_29),
  .I0(mux_o_26),
  .I1(mux_o_27),
  .S0(rad[7])
);
MUX2 mux_inst_30 (
  .O(dout[0]),
  .I0(mux_o_28),
  .I1(mux_o_29),
  .S0(rad[8])
);
MUX2 mux_inst_31 (
  .O(mux_o_31),
  .I0(ram16sdp_inst_0_dout[1]),
  .I1(ram16sdp_inst_2_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_32 (
  .O(mux_o_32),
  .I0(ram16sdp_inst_4_dout[1]),
  .I1(ram16sdp_inst_6_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_33 (
  .O(mux_o_33),
  .I0(ram16sdp_inst_8_dout[1]),
  .I1(ram16sdp_inst_10_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_34 (
  .O(mux_o_34),
  .I0(ram16sdp_inst_12_dout[1]),
  .I1(ram16sdp_inst_14_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_35 (
  .O(mux_o_35),
  .I0(ram16sdp_inst_16_dout[1]),
  .I1(ram16sdp_inst_18_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_36 (
  .O(mux_o_36),
  .I0(ram16sdp_inst_20_dout[1]),
  .I1(ram16sdp_inst_22_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_37 (
  .O(mux_o_37),
  .I0(ram16sdp_inst_24_dout[1]),
  .I1(ram16sdp_inst_26_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_38 (
  .O(mux_o_38),
  .I0(ram16sdp_inst_28_dout[1]),
  .I1(ram16sdp_inst_30_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_39 (
  .O(mux_o_39),
  .I0(ram16sdp_inst_32_dout[1]),
  .I1(ram16sdp_inst_34_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_40 (
  .O(mux_o_40),
  .I0(ram16sdp_inst_36_dout[1]),
  .I1(ram16sdp_inst_38_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_41 (
  .O(mux_o_41),
  .I0(ram16sdp_inst_40_dout[1]),
  .I1(ram16sdp_inst_42_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_42 (
  .O(mux_o_42),
  .I0(ram16sdp_inst_44_dout[1]),
  .I1(ram16sdp_inst_46_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_43 (
  .O(mux_o_43),
  .I0(ram16sdp_inst_48_dout[1]),
  .I1(ram16sdp_inst_50_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_44 (
  .O(mux_o_44),
  .I0(ram16sdp_inst_52_dout[1]),
  .I1(ram16sdp_inst_54_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_45 (
  .O(mux_o_45),
  .I0(ram16sdp_inst_56_dout[1]),
  .I1(ram16sdp_inst_58_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_46 (
  .O(mux_o_46),
  .I0(ram16sdp_inst_60_dout[1]),
  .I1(ram16sdp_inst_62_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_47 (
  .O(mux_o_47),
  .I0(mux_o_31),
  .I1(mux_o_32),
  .S0(rad[5])
);
MUX2 mux_inst_48 (
  .O(mux_o_48),
  .I0(mux_o_33),
  .I1(mux_o_34),
  .S0(rad[5])
);
MUX2 mux_inst_49 (
  .O(mux_o_49),
  .I0(mux_o_35),
  .I1(mux_o_36),
  .S0(rad[5])
);
MUX2 mux_inst_50 (
  .O(mux_o_50),
  .I0(mux_o_37),
  .I1(mux_o_38),
  .S0(rad[5])
);
MUX2 mux_inst_51 (
  .O(mux_o_51),
  .I0(mux_o_39),
  .I1(mux_o_40),
  .S0(rad[5])
);
MUX2 mux_inst_52 (
  .O(mux_o_52),
  .I0(mux_o_41),
  .I1(mux_o_42),
  .S0(rad[5])
);
MUX2 mux_inst_53 (
  .O(mux_o_53),
  .I0(mux_o_43),
  .I1(mux_o_44),
  .S0(rad[5])
);
MUX2 mux_inst_54 (
  .O(mux_o_54),
  .I0(mux_o_45),
  .I1(mux_o_46),
  .S0(rad[5])
);
MUX2 mux_inst_55 (
  .O(mux_o_55),
  .I0(mux_o_47),
  .I1(mux_o_48),
  .S0(rad[6])
);
MUX2 mux_inst_56 (
  .O(mux_o_56),
  .I0(mux_o_49),
  .I1(mux_o_50),
  .S0(rad[6])
);
MUX2 mux_inst_57 (
  .O(mux_o_57),
  .I0(mux_o_51),
  .I1(mux_o_52),
  .S0(rad[6])
);
MUX2 mux_inst_58 (
  .O(mux_o_58),
  .I0(mux_o_53),
  .I1(mux_o_54),
  .S0(rad[6])
);
MUX2 mux_inst_59 (
  .O(mux_o_59),
  .I0(mux_o_55),
  .I1(mux_o_56),
  .S0(rad[7])
);
MUX2 mux_inst_60 (
  .O(mux_o_60),
  .I0(mux_o_57),
  .I1(mux_o_58),
  .S0(rad[7])
);
MUX2 mux_inst_61 (
  .O(dout[1]),
  .I0(mux_o_59),
  .I1(mux_o_60),
  .S0(rad[8])
);
MUX2 mux_inst_62 (
  .O(mux_o_62),
  .I0(ram16sdp_inst_0_dout[2]),
  .I1(ram16sdp_inst_2_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_63 (
  .O(mux_o_63),
  .I0(ram16sdp_inst_4_dout[2]),
  .I1(ram16sdp_inst_6_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_64 (
  .O(mux_o_64),
  .I0(ram16sdp_inst_8_dout[2]),
  .I1(ram16sdp_inst_10_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_65 (
  .O(mux_o_65),
  .I0(ram16sdp_inst_12_dout[2]),
  .I1(ram16sdp_inst_14_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_66 (
  .O(mux_o_66),
  .I0(ram16sdp_inst_16_dout[2]),
  .I1(ram16sdp_inst_18_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_67 (
  .O(mux_o_67),
  .I0(ram16sdp_inst_20_dout[2]),
  .I1(ram16sdp_inst_22_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_68 (
  .O(mux_o_68),
  .I0(ram16sdp_inst_24_dout[2]),
  .I1(ram16sdp_inst_26_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_69 (
  .O(mux_o_69),
  .I0(ram16sdp_inst_28_dout[2]),
  .I1(ram16sdp_inst_30_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_70 (
  .O(mux_o_70),
  .I0(ram16sdp_inst_32_dout[2]),
  .I1(ram16sdp_inst_34_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_71 (
  .O(mux_o_71),
  .I0(ram16sdp_inst_36_dout[2]),
  .I1(ram16sdp_inst_38_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_72 (
  .O(mux_o_72),
  .I0(ram16sdp_inst_40_dout[2]),
  .I1(ram16sdp_inst_42_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_73 (
  .O(mux_o_73),
  .I0(ram16sdp_inst_44_dout[2]),
  .I1(ram16sdp_inst_46_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_74 (
  .O(mux_o_74),
  .I0(ram16sdp_inst_48_dout[2]),
  .I1(ram16sdp_inst_50_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_75 (
  .O(mux_o_75),
  .I0(ram16sdp_inst_52_dout[2]),
  .I1(ram16sdp_inst_54_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_76 (
  .O(mux_o_76),
  .I0(ram16sdp_inst_56_dout[2]),
  .I1(ram16sdp_inst_58_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_77 (
  .O(mux_o_77),
  .I0(ram16sdp_inst_60_dout[2]),
  .I1(ram16sdp_inst_62_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_78 (
  .O(mux_o_78),
  .I0(mux_o_62),
  .I1(mux_o_63),
  .S0(rad[5])
);
MUX2 mux_inst_79 (
  .O(mux_o_79),
  .I0(mux_o_64),
  .I1(mux_o_65),
  .S0(rad[5])
);
MUX2 mux_inst_80 (
  .O(mux_o_80),
  .I0(mux_o_66),
  .I1(mux_o_67),
  .S0(rad[5])
);
MUX2 mux_inst_81 (
  .O(mux_o_81),
  .I0(mux_o_68),
  .I1(mux_o_69),
  .S0(rad[5])
);
MUX2 mux_inst_82 (
  .O(mux_o_82),
  .I0(mux_o_70),
  .I1(mux_o_71),
  .S0(rad[5])
);
MUX2 mux_inst_83 (
  .O(mux_o_83),
  .I0(mux_o_72),
  .I1(mux_o_73),
  .S0(rad[5])
);
MUX2 mux_inst_84 (
  .O(mux_o_84),
  .I0(mux_o_74),
  .I1(mux_o_75),
  .S0(rad[5])
);
MUX2 mux_inst_85 (
  .O(mux_o_85),
  .I0(mux_o_76),
  .I1(mux_o_77),
  .S0(rad[5])
);
MUX2 mux_inst_86 (
  .O(mux_o_86),
  .I0(mux_o_78),
  .I1(mux_o_79),
  .S0(rad[6])
);
MUX2 mux_inst_87 (
  .O(mux_o_87),
  .I0(mux_o_80),
  .I1(mux_o_81),
  .S0(rad[6])
);
MUX2 mux_inst_88 (
  .O(mux_o_88),
  .I0(mux_o_82),
  .I1(mux_o_83),
  .S0(rad[6])
);
MUX2 mux_inst_89 (
  .O(mux_o_89),
  .I0(mux_o_84),
  .I1(mux_o_85),
  .S0(rad[6])
);
MUX2 mux_inst_90 (
  .O(mux_o_90),
  .I0(mux_o_86),
  .I1(mux_o_87),
  .S0(rad[7])
);
MUX2 mux_inst_91 (
  .O(mux_o_91),
  .I0(mux_o_88),
  .I1(mux_o_89),
  .S0(rad[7])
);
MUX2 mux_inst_92 (
  .O(dout[2]),
  .I0(mux_o_90),
  .I1(mux_o_91),
  .S0(rad[8])
);
MUX2 mux_inst_93 (
  .O(mux_o_93),
  .I0(ram16sdp_inst_0_dout[3]),
  .I1(ram16sdp_inst_2_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_94 (
  .O(mux_o_94),
  .I0(ram16sdp_inst_4_dout[3]),
  .I1(ram16sdp_inst_6_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_95 (
  .O(mux_o_95),
  .I0(ram16sdp_inst_8_dout[3]),
  .I1(ram16sdp_inst_10_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_96 (
  .O(mux_o_96),
  .I0(ram16sdp_inst_12_dout[3]),
  .I1(ram16sdp_inst_14_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_97 (
  .O(mux_o_97),
  .I0(ram16sdp_inst_16_dout[3]),
  .I1(ram16sdp_inst_18_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_98 (
  .O(mux_o_98),
  .I0(ram16sdp_inst_20_dout[3]),
  .I1(ram16sdp_inst_22_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_99 (
  .O(mux_o_99),
  .I0(ram16sdp_inst_24_dout[3]),
  .I1(ram16sdp_inst_26_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_100 (
  .O(mux_o_100),
  .I0(ram16sdp_inst_28_dout[3]),
  .I1(ram16sdp_inst_30_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_101 (
  .O(mux_o_101),
  .I0(ram16sdp_inst_32_dout[3]),
  .I1(ram16sdp_inst_34_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_102 (
  .O(mux_o_102),
  .I0(ram16sdp_inst_36_dout[3]),
  .I1(ram16sdp_inst_38_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_103 (
  .O(mux_o_103),
  .I0(ram16sdp_inst_40_dout[3]),
  .I1(ram16sdp_inst_42_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_104 (
  .O(mux_o_104),
  .I0(ram16sdp_inst_44_dout[3]),
  .I1(ram16sdp_inst_46_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_105 (
  .O(mux_o_105),
  .I0(ram16sdp_inst_48_dout[3]),
  .I1(ram16sdp_inst_50_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_106 (
  .O(mux_o_106),
  .I0(ram16sdp_inst_52_dout[3]),
  .I1(ram16sdp_inst_54_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_107 (
  .O(mux_o_107),
  .I0(ram16sdp_inst_56_dout[3]),
  .I1(ram16sdp_inst_58_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_108 (
  .O(mux_o_108),
  .I0(ram16sdp_inst_60_dout[3]),
  .I1(ram16sdp_inst_62_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_109 (
  .O(mux_o_109),
  .I0(mux_o_93),
  .I1(mux_o_94),
  .S0(rad[5])
);
MUX2 mux_inst_110 (
  .O(mux_o_110),
  .I0(mux_o_95),
  .I1(mux_o_96),
  .S0(rad[5])
);
MUX2 mux_inst_111 (
  .O(mux_o_111),
  .I0(mux_o_97),
  .I1(mux_o_98),
  .S0(rad[5])
);
MUX2 mux_inst_112 (
  .O(mux_o_112),
  .I0(mux_o_99),
  .I1(mux_o_100),
  .S0(rad[5])
);
MUX2 mux_inst_113 (
  .O(mux_o_113),
  .I0(mux_o_101),
  .I1(mux_o_102),
  .S0(rad[5])
);
MUX2 mux_inst_114 (
  .O(mux_o_114),
  .I0(mux_o_103),
  .I1(mux_o_104),
  .S0(rad[5])
);
MUX2 mux_inst_115 (
  .O(mux_o_115),
  .I0(mux_o_105),
  .I1(mux_o_106),
  .S0(rad[5])
);
MUX2 mux_inst_116 (
  .O(mux_o_116),
  .I0(mux_o_107),
  .I1(mux_o_108),
  .S0(rad[5])
);
MUX2 mux_inst_117 (
  .O(mux_o_117),
  .I0(mux_o_109),
  .I1(mux_o_110),
  .S0(rad[6])
);
MUX2 mux_inst_118 (
  .O(mux_o_118),
  .I0(mux_o_111),
  .I1(mux_o_112),
  .S0(rad[6])
);
MUX2 mux_inst_119 (
  .O(mux_o_119),
  .I0(mux_o_113),
  .I1(mux_o_114),
  .S0(rad[6])
);
MUX2 mux_inst_120 (
  .O(mux_o_120),
  .I0(mux_o_115),
  .I1(mux_o_116),
  .S0(rad[6])
);
MUX2 mux_inst_121 (
  .O(mux_o_121),
  .I0(mux_o_117),
  .I1(mux_o_118),
  .S0(rad[7])
);
MUX2 mux_inst_122 (
  .O(mux_o_122),
  .I0(mux_o_119),
  .I1(mux_o_120),
  .S0(rad[7])
);
MUX2 mux_inst_123 (
  .O(dout[3]),
  .I0(mux_o_121),
  .I1(mux_o_122),
  .S0(rad[8])
);
MUX2 mux_inst_124 (
  .O(mux_o_124),
  .I0(ram16sdp_inst_1_dout[4]),
  .I1(ram16sdp_inst_3_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_125 (
  .O(mux_o_125),
  .I0(ram16sdp_inst_5_dout[4]),
  .I1(ram16sdp_inst_7_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_126 (
  .O(mux_o_126),
  .I0(ram16sdp_inst_9_dout[4]),
  .I1(ram16sdp_inst_11_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_127 (
  .O(mux_o_127),
  .I0(ram16sdp_inst_13_dout[4]),
  .I1(ram16sdp_inst_15_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_128 (
  .O(mux_o_128),
  .I0(ram16sdp_inst_17_dout[4]),
  .I1(ram16sdp_inst_19_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_129 (
  .O(mux_o_129),
  .I0(ram16sdp_inst_21_dout[4]),
  .I1(ram16sdp_inst_23_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_130 (
  .O(mux_o_130),
  .I0(ram16sdp_inst_25_dout[4]),
  .I1(ram16sdp_inst_27_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_131 (
  .O(mux_o_131),
  .I0(ram16sdp_inst_29_dout[4]),
  .I1(ram16sdp_inst_31_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_132 (
  .O(mux_o_132),
  .I0(ram16sdp_inst_33_dout[4]),
  .I1(ram16sdp_inst_35_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_133 (
  .O(mux_o_133),
  .I0(ram16sdp_inst_37_dout[4]),
  .I1(ram16sdp_inst_39_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_134 (
  .O(mux_o_134),
  .I0(ram16sdp_inst_41_dout[4]),
  .I1(ram16sdp_inst_43_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_135 (
  .O(mux_o_135),
  .I0(ram16sdp_inst_45_dout[4]),
  .I1(ram16sdp_inst_47_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_136 (
  .O(mux_o_136),
  .I0(ram16sdp_inst_49_dout[4]),
  .I1(ram16sdp_inst_51_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_137 (
  .O(mux_o_137),
  .I0(ram16sdp_inst_53_dout[4]),
  .I1(ram16sdp_inst_55_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_138 (
  .O(mux_o_138),
  .I0(ram16sdp_inst_57_dout[4]),
  .I1(ram16sdp_inst_59_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_139 (
  .O(mux_o_139),
  .I0(ram16sdp_inst_61_dout[4]),
  .I1(ram16sdp_inst_63_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_140 (
  .O(mux_o_140),
  .I0(mux_o_124),
  .I1(mux_o_125),
  .S0(rad[5])
);
MUX2 mux_inst_141 (
  .O(mux_o_141),
  .I0(mux_o_126),
  .I1(mux_o_127),
  .S0(rad[5])
);
MUX2 mux_inst_142 (
  .O(mux_o_142),
  .I0(mux_o_128),
  .I1(mux_o_129),
  .S0(rad[5])
);
MUX2 mux_inst_143 (
  .O(mux_o_143),
  .I0(mux_o_130),
  .I1(mux_o_131),
  .S0(rad[5])
);
MUX2 mux_inst_144 (
  .O(mux_o_144),
  .I0(mux_o_132),
  .I1(mux_o_133),
  .S0(rad[5])
);
MUX2 mux_inst_145 (
  .O(mux_o_145),
  .I0(mux_o_134),
  .I1(mux_o_135),
  .S0(rad[5])
);
MUX2 mux_inst_146 (
  .O(mux_o_146),
  .I0(mux_o_136),
  .I1(mux_o_137),
  .S0(rad[5])
);
MUX2 mux_inst_147 (
  .O(mux_o_147),
  .I0(mux_o_138),
  .I1(mux_o_139),
  .S0(rad[5])
);
MUX2 mux_inst_148 (
  .O(mux_o_148),
  .I0(mux_o_140),
  .I1(mux_o_141),
  .S0(rad[6])
);
MUX2 mux_inst_149 (
  .O(mux_o_149),
  .I0(mux_o_142),
  .I1(mux_o_143),
  .S0(rad[6])
);
MUX2 mux_inst_150 (
  .O(mux_o_150),
  .I0(mux_o_144),
  .I1(mux_o_145),
  .S0(rad[6])
);
MUX2 mux_inst_151 (
  .O(mux_o_151),
  .I0(mux_o_146),
  .I1(mux_o_147),
  .S0(rad[6])
);
MUX2 mux_inst_152 (
  .O(mux_o_152),
  .I0(mux_o_148),
  .I1(mux_o_149),
  .S0(rad[7])
);
MUX2 mux_inst_153 (
  .O(mux_o_153),
  .I0(mux_o_150),
  .I1(mux_o_151),
  .S0(rad[7])
);
MUX2 mux_inst_154 (
  .O(dout[4]),
  .I0(mux_o_152),
  .I1(mux_o_153),
  .S0(rad[8])
);
MUX2 mux_inst_155 (
  .O(mux_o_155),
  .I0(ram16sdp_inst_1_dout[5]),
  .I1(ram16sdp_inst_3_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_156 (
  .O(mux_o_156),
  .I0(ram16sdp_inst_5_dout[5]),
  .I1(ram16sdp_inst_7_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_157 (
  .O(mux_o_157),
  .I0(ram16sdp_inst_9_dout[5]),
  .I1(ram16sdp_inst_11_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_158 (
  .O(mux_o_158),
  .I0(ram16sdp_inst_13_dout[5]),
  .I1(ram16sdp_inst_15_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_159 (
  .O(mux_o_159),
  .I0(ram16sdp_inst_17_dout[5]),
  .I1(ram16sdp_inst_19_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_160 (
  .O(mux_o_160),
  .I0(ram16sdp_inst_21_dout[5]),
  .I1(ram16sdp_inst_23_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_161 (
  .O(mux_o_161),
  .I0(ram16sdp_inst_25_dout[5]),
  .I1(ram16sdp_inst_27_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_162 (
  .O(mux_o_162),
  .I0(ram16sdp_inst_29_dout[5]),
  .I1(ram16sdp_inst_31_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_163 (
  .O(mux_o_163),
  .I0(ram16sdp_inst_33_dout[5]),
  .I1(ram16sdp_inst_35_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_164 (
  .O(mux_o_164),
  .I0(ram16sdp_inst_37_dout[5]),
  .I1(ram16sdp_inst_39_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_165 (
  .O(mux_o_165),
  .I0(ram16sdp_inst_41_dout[5]),
  .I1(ram16sdp_inst_43_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_166 (
  .O(mux_o_166),
  .I0(ram16sdp_inst_45_dout[5]),
  .I1(ram16sdp_inst_47_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_167 (
  .O(mux_o_167),
  .I0(ram16sdp_inst_49_dout[5]),
  .I1(ram16sdp_inst_51_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_168 (
  .O(mux_o_168),
  .I0(ram16sdp_inst_53_dout[5]),
  .I1(ram16sdp_inst_55_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_169 (
  .O(mux_o_169),
  .I0(ram16sdp_inst_57_dout[5]),
  .I1(ram16sdp_inst_59_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_170 (
  .O(mux_o_170),
  .I0(ram16sdp_inst_61_dout[5]),
  .I1(ram16sdp_inst_63_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_171 (
  .O(mux_o_171),
  .I0(mux_o_155),
  .I1(mux_o_156),
  .S0(rad[5])
);
MUX2 mux_inst_172 (
  .O(mux_o_172),
  .I0(mux_o_157),
  .I1(mux_o_158),
  .S0(rad[5])
);
MUX2 mux_inst_173 (
  .O(mux_o_173),
  .I0(mux_o_159),
  .I1(mux_o_160),
  .S0(rad[5])
);
MUX2 mux_inst_174 (
  .O(mux_o_174),
  .I0(mux_o_161),
  .I1(mux_o_162),
  .S0(rad[5])
);
MUX2 mux_inst_175 (
  .O(mux_o_175),
  .I0(mux_o_163),
  .I1(mux_o_164),
  .S0(rad[5])
);
MUX2 mux_inst_176 (
  .O(mux_o_176),
  .I0(mux_o_165),
  .I1(mux_o_166),
  .S0(rad[5])
);
MUX2 mux_inst_177 (
  .O(mux_o_177),
  .I0(mux_o_167),
  .I1(mux_o_168),
  .S0(rad[5])
);
MUX2 mux_inst_178 (
  .O(mux_o_178),
  .I0(mux_o_169),
  .I1(mux_o_170),
  .S0(rad[5])
);
MUX2 mux_inst_179 (
  .O(mux_o_179),
  .I0(mux_o_171),
  .I1(mux_o_172),
  .S0(rad[6])
);
MUX2 mux_inst_180 (
  .O(mux_o_180),
  .I0(mux_o_173),
  .I1(mux_o_174),
  .S0(rad[6])
);
MUX2 mux_inst_181 (
  .O(mux_o_181),
  .I0(mux_o_175),
  .I1(mux_o_176),
  .S0(rad[6])
);
MUX2 mux_inst_182 (
  .O(mux_o_182),
  .I0(mux_o_177),
  .I1(mux_o_178),
  .S0(rad[6])
);
MUX2 mux_inst_183 (
  .O(mux_o_183),
  .I0(mux_o_179),
  .I1(mux_o_180),
  .S0(rad[7])
);
MUX2 mux_inst_184 (
  .O(mux_o_184),
  .I0(mux_o_181),
  .I1(mux_o_182),
  .S0(rad[7])
);
MUX2 mux_inst_185 (
  .O(dout[5]),
  .I0(mux_o_183),
  .I1(mux_o_184),
  .S0(rad[8])
);
MUX2 mux_inst_186 (
  .O(mux_o_186),
  .I0(ram16sdp_inst_1_dout[6]),
  .I1(ram16sdp_inst_3_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_187 (
  .O(mux_o_187),
  .I0(ram16sdp_inst_5_dout[6]),
  .I1(ram16sdp_inst_7_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_188 (
  .O(mux_o_188),
  .I0(ram16sdp_inst_9_dout[6]),
  .I1(ram16sdp_inst_11_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_189 (
  .O(mux_o_189),
  .I0(ram16sdp_inst_13_dout[6]),
  .I1(ram16sdp_inst_15_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_190 (
  .O(mux_o_190),
  .I0(ram16sdp_inst_17_dout[6]),
  .I1(ram16sdp_inst_19_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_191 (
  .O(mux_o_191),
  .I0(ram16sdp_inst_21_dout[6]),
  .I1(ram16sdp_inst_23_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_192 (
  .O(mux_o_192),
  .I0(ram16sdp_inst_25_dout[6]),
  .I1(ram16sdp_inst_27_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_193 (
  .O(mux_o_193),
  .I0(ram16sdp_inst_29_dout[6]),
  .I1(ram16sdp_inst_31_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_194 (
  .O(mux_o_194),
  .I0(ram16sdp_inst_33_dout[6]),
  .I1(ram16sdp_inst_35_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_195 (
  .O(mux_o_195),
  .I0(ram16sdp_inst_37_dout[6]),
  .I1(ram16sdp_inst_39_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_196 (
  .O(mux_o_196),
  .I0(ram16sdp_inst_41_dout[6]),
  .I1(ram16sdp_inst_43_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_197 (
  .O(mux_o_197),
  .I0(ram16sdp_inst_45_dout[6]),
  .I1(ram16sdp_inst_47_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_198 (
  .O(mux_o_198),
  .I0(ram16sdp_inst_49_dout[6]),
  .I1(ram16sdp_inst_51_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_199 (
  .O(mux_o_199),
  .I0(ram16sdp_inst_53_dout[6]),
  .I1(ram16sdp_inst_55_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_200 (
  .O(mux_o_200),
  .I0(ram16sdp_inst_57_dout[6]),
  .I1(ram16sdp_inst_59_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_201 (
  .O(mux_o_201),
  .I0(ram16sdp_inst_61_dout[6]),
  .I1(ram16sdp_inst_63_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_202 (
  .O(mux_o_202),
  .I0(mux_o_186),
  .I1(mux_o_187),
  .S0(rad[5])
);
MUX2 mux_inst_203 (
  .O(mux_o_203),
  .I0(mux_o_188),
  .I1(mux_o_189),
  .S0(rad[5])
);
MUX2 mux_inst_204 (
  .O(mux_o_204),
  .I0(mux_o_190),
  .I1(mux_o_191),
  .S0(rad[5])
);
MUX2 mux_inst_205 (
  .O(mux_o_205),
  .I0(mux_o_192),
  .I1(mux_o_193),
  .S0(rad[5])
);
MUX2 mux_inst_206 (
  .O(mux_o_206),
  .I0(mux_o_194),
  .I1(mux_o_195),
  .S0(rad[5])
);
MUX2 mux_inst_207 (
  .O(mux_o_207),
  .I0(mux_o_196),
  .I1(mux_o_197),
  .S0(rad[5])
);
MUX2 mux_inst_208 (
  .O(mux_o_208),
  .I0(mux_o_198),
  .I1(mux_o_199),
  .S0(rad[5])
);
MUX2 mux_inst_209 (
  .O(mux_o_209),
  .I0(mux_o_200),
  .I1(mux_o_201),
  .S0(rad[5])
);
MUX2 mux_inst_210 (
  .O(mux_o_210),
  .I0(mux_o_202),
  .I1(mux_o_203),
  .S0(rad[6])
);
MUX2 mux_inst_211 (
  .O(mux_o_211),
  .I0(mux_o_204),
  .I1(mux_o_205),
  .S0(rad[6])
);
MUX2 mux_inst_212 (
  .O(mux_o_212),
  .I0(mux_o_206),
  .I1(mux_o_207),
  .S0(rad[6])
);
MUX2 mux_inst_213 (
  .O(mux_o_213),
  .I0(mux_o_208),
  .I1(mux_o_209),
  .S0(rad[6])
);
MUX2 mux_inst_214 (
  .O(mux_o_214),
  .I0(mux_o_210),
  .I1(mux_o_211),
  .S0(rad[7])
);
MUX2 mux_inst_215 (
  .O(mux_o_215),
  .I0(mux_o_212),
  .I1(mux_o_213),
  .S0(rad[7])
);
MUX2 mux_inst_216 (
  .O(dout[6]),
  .I0(mux_o_214),
  .I1(mux_o_215),
  .S0(rad[8])
);
MUX2 mux_inst_217 (
  .O(mux_o_217),
  .I0(ram16sdp_inst_1_dout[7]),
  .I1(ram16sdp_inst_3_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_218 (
  .O(mux_o_218),
  .I0(ram16sdp_inst_5_dout[7]),
  .I1(ram16sdp_inst_7_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_219 (
  .O(mux_o_219),
  .I0(ram16sdp_inst_9_dout[7]),
  .I1(ram16sdp_inst_11_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_220 (
  .O(mux_o_220),
  .I0(ram16sdp_inst_13_dout[7]),
  .I1(ram16sdp_inst_15_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_221 (
  .O(mux_o_221),
  .I0(ram16sdp_inst_17_dout[7]),
  .I1(ram16sdp_inst_19_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_222 (
  .O(mux_o_222),
  .I0(ram16sdp_inst_21_dout[7]),
  .I1(ram16sdp_inst_23_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_223 (
  .O(mux_o_223),
  .I0(ram16sdp_inst_25_dout[7]),
  .I1(ram16sdp_inst_27_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_224 (
  .O(mux_o_224),
  .I0(ram16sdp_inst_29_dout[7]),
  .I1(ram16sdp_inst_31_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_225 (
  .O(mux_o_225),
  .I0(ram16sdp_inst_33_dout[7]),
  .I1(ram16sdp_inst_35_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_226 (
  .O(mux_o_226),
  .I0(ram16sdp_inst_37_dout[7]),
  .I1(ram16sdp_inst_39_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_227 (
  .O(mux_o_227),
  .I0(ram16sdp_inst_41_dout[7]),
  .I1(ram16sdp_inst_43_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_228 (
  .O(mux_o_228),
  .I0(ram16sdp_inst_45_dout[7]),
  .I1(ram16sdp_inst_47_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_229 (
  .O(mux_o_229),
  .I0(ram16sdp_inst_49_dout[7]),
  .I1(ram16sdp_inst_51_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_230 (
  .O(mux_o_230),
  .I0(ram16sdp_inst_53_dout[7]),
  .I1(ram16sdp_inst_55_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_231 (
  .O(mux_o_231),
  .I0(ram16sdp_inst_57_dout[7]),
  .I1(ram16sdp_inst_59_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_232 (
  .O(mux_o_232),
  .I0(ram16sdp_inst_61_dout[7]),
  .I1(ram16sdp_inst_63_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_233 (
  .O(mux_o_233),
  .I0(mux_o_217),
  .I1(mux_o_218),
  .S0(rad[5])
);
MUX2 mux_inst_234 (
  .O(mux_o_234),
  .I0(mux_o_219),
  .I1(mux_o_220),
  .S0(rad[5])
);
MUX2 mux_inst_235 (
  .O(mux_o_235),
  .I0(mux_o_221),
  .I1(mux_o_222),
  .S0(rad[5])
);
MUX2 mux_inst_236 (
  .O(mux_o_236),
  .I0(mux_o_223),
  .I1(mux_o_224),
  .S0(rad[5])
);
MUX2 mux_inst_237 (
  .O(mux_o_237),
  .I0(mux_o_225),
  .I1(mux_o_226),
  .S0(rad[5])
);
MUX2 mux_inst_238 (
  .O(mux_o_238),
  .I0(mux_o_227),
  .I1(mux_o_228),
  .S0(rad[5])
);
MUX2 mux_inst_239 (
  .O(mux_o_239),
  .I0(mux_o_229),
  .I1(mux_o_230),
  .S0(rad[5])
);
MUX2 mux_inst_240 (
  .O(mux_o_240),
  .I0(mux_o_231),
  .I1(mux_o_232),
  .S0(rad[5])
);
MUX2 mux_inst_241 (
  .O(mux_o_241),
  .I0(mux_o_233),
  .I1(mux_o_234),
  .S0(rad[6])
);
MUX2 mux_inst_242 (
  .O(mux_o_242),
  .I0(mux_o_235),
  .I1(mux_o_236),
  .S0(rad[6])
);
MUX2 mux_inst_243 (
  .O(mux_o_243),
  .I0(mux_o_237),
  .I1(mux_o_238),
  .S0(rad[6])
);
MUX2 mux_inst_244 (
  .O(mux_o_244),
  .I0(mux_o_239),
  .I1(mux_o_240),
  .S0(rad[6])
);
MUX2 mux_inst_245 (
  .O(mux_o_245),
  .I0(mux_o_241),
  .I1(mux_o_242),
  .S0(rad[7])
);
MUX2 mux_inst_246 (
  .O(mux_o_246),
  .I0(mux_o_243),
  .I1(mux_o_244),
  .S0(rad[7])
);
MUX2 mux_inst_247 (
  .O(dout[7]),
  .I0(mux_o_245),
  .I1(mux_o_246),
  .S0(rad[8])
);
endmodule //usb_retrans_ram
