`define MODULE_NAME mult_signed_nuc
`define SIGNED_A
`define SIGNED_B
`define DATA_B
`define LUT
`define PIPELINE
